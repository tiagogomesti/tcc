----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:59:18 02/18/2015 
-- Design Name: 
-- Module Name:    command_tb - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.toneDetectorPackage.all;



entity command_tb is
port
(
	RESET								: in std_logic;
	CLK									: in std_logic;

	CMD_TX_DATA					: out unsigned (WORD_SIZE-1 downto 0);
	CMD_WORD_INDEX			: out integer range 0 to 6;
	WRITE_CMD_BUFFER	: out	std_logic;
	CMD_TX							: out std_logic;
	CMD_TX_ACK					: in std_logic
);

end command_tb;

architecture Behavioral of command_tb is

begin


	process
	begin
		wait until RESET = '0';

		CMD_TX <= '1'; 

		wait until CMD_TX_ACK = '1';

		wait for CLOCK_PERIOD;

		CMD_WORD_INDEX <= 0;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"0001";
		WRITE_CMD_BUFFER <= '1';

		CMD_WORD_INDEX <= 1;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"0025";

		CMD_WORD_INDEX <= 2;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"0000";

		CMD_WORD_INDEX <= 3;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"0300";

		CMD_WORD_INDEX <= 4;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"0015";

		CMD_WORD_INDEX <= 5;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"7942";

		CMD_WORD_INDEX <= 6;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"789a";

		wait for CLOCK_PERIOD;

		WRITE_CMD_BUFFER <= '0';
		CMD_TX <= '0';


		wait for CLOCK_PERIOD;

		wait for CLOCK_PERIOD;

		wait for CLOCK_PERIOD;


--=======================================--
		CMD_TX <= '1'; 

		wait until CMD_TX_ACK = '1';

		wait for CLOCK_PERIOD;

		CMD_WORD_INDEX <= 0;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"0003";
		WRITE_CMD_BUFFER <= '1';

		CMD_WORD_INDEX <= 1;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"0025";

		CMD_WORD_INDEX <= 2;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"0000";

		CMD_WORD_INDEX <= 3;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"0300";

		CMD_WORD_INDEX <= 4;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"0015";

		CMD_WORD_INDEX <= 5;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"7942";

		CMD_WORD_INDEX <= 6;
		wait for CLOCK_PERIOD;
		CMD_TX_DATA	<= x"789a";

		CMD_TX <= '0';



		wait;


	end process;



end Behavioral;

